//Simple verilod display module.

module disp();
	initial
	$display("Verilog Display");
endmodule
